library verilog;
use verilog.vl_types.all;
entity contador_p3_vlg_sample_tst is
    port(
        clock           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end contador_p3_vlg_sample_tst;
