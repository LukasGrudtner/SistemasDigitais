library verilog;
use verilog.vl_types.all;
entity part5_vlg_vec_tst is
end part5_vlg_vec_tst;
